module main(CLK,TXD,RXD,LED);
	input CLK;
	input TXD;
	output RXD;
	output LED;
endmodule
